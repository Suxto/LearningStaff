library verilog;
use verilog.vl_types.all;
entity TestRam_vlg_check_tst is
    port(
        DBus            : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end TestRam_vlg_check_tst;
