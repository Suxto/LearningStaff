library verilog;
use verilog.vl_types.all;
entity Calc_vlg_vec_tst is
end Calc_vlg_vec_tst;
