library verilog;
use verilog.vl_types.all;
entity StaticLED_vlg_vec_tst is
end StaticLED_vlg_vec_tst;
