library verilog;
use verilog.vl_types.all;
entity register_led_vlg_vec_tst is
end register_led_vlg_vec_tst;
