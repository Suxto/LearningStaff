library verilog;
use verilog.vl_types.all;
entity mux4_vlg_vec_tst is
end mux4_vlg_vec_tst;
