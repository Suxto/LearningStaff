library verilog;
use verilog.vl_types.all;
entity TestRam_vlg_vec_tst is
end TestRam_vlg_vec_tst;
