library verilog;
use verilog.vl_types.all;
entity Time_vlg_vec_tst is
end Time_vlg_vec_tst;
