library verilog;
use verilog.vl_types.all;
entity latch_8bit_vlg_vec_tst is
end latch_8bit_vlg_vec_tst;
