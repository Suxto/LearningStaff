library verilog;
use verilog.vl_types.all;
entity mux8_vlg_vec_tst is
end mux8_vlg_vec_tst;
